`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.02.2024 11:55:31
// Design Name: 
// Module Name: bram
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module bram	#(
	parameter WIDTH = 32,
	parameter DEPTH  = 10,
	parameter MEM_READ_PORTS = 2
	) (
		input clk,                                        // Señal de reloj
		input rst,                                        // Señal de reset
		input [(DEPTH*MEM_READ_PORTS)-1:0] addr_read,     // Dirección de lectura (anchura varia segun numero de puertos de lectura)
		input [DEPTH-1:0] addr_write,                     // Direccion de escritura
		input [WIDTH-1:0] data,                           // Dato entrante de escritura
		input w_en,                                       // Señal de escritura
		output [(WIDTH*MEM_READ_PORTS)-1:0] rd_o          // Salida de datos (anchura varia segun numero de puertos de lectura)
    );
    
    reg [WIDTH-1:0] mem [0:2**DEPTH-1];     // Memoria
    
    // Bloque always para gestionar la escritura de memoria
    // Señal de reset -> se reinicia el contenido a 0 (y se escriben algunos datos usados para pruebas)
    // Señal de escritura -> se escribe el dato entrante "data" en la posición apuntada por addr_write
    integer rst_mem;
    always @(posedge clk) begin
    	if (rst) begin
    		for(rst_mem = 0; rst_mem < 2**DEPTH; rst_mem = rst_mem + 1) begin
    			mem[rst_mem] <= 0;
    		end
			mem[0] <=   32'b00111111100000000000000000000000;    //   1;
			mem[1] <=   32'b01000000100000000000000000000000;    //   4;  
			mem[2] <=   32'b01000001000100000000000000000000;    //   9;
			mem[3] <=   32'b01000001100000000000000000000000;    //  16;
			mem[4] <=   32'b01000001110010000000000000000000;    //  25;
			mem[5] <=   32'b01000010000100000000000000000000;    //  36;
			mem[6] <=   32'b01000010010001000000000000000000;    //  49;
			mem[7] <=   32'b01000010100000000000000000000000;    //  64;    /* 32'b10000000000000000000000000000000; */
			mem[8] <=   32'b0_00000000_00000000000000000000000;  // 2;
			mem[9] <=   32'b0_10000000_00000000000000000000000;  // 4;
			mem[10] <=  32'b0_00000000_00000000000000000000000;  // 2;
			mem[11] <=  32'b0_10000000_00000000000000000000000;  // 2;
			mem[12] <=  32'b0_00000000_00000000000000000000000;  // 2;
			mem[13] <=  32'b0_10000000_00000000000000000000000;  // 2;
			mem[14] <=  32'b0_00000000_00000000000000000000000;  // 2;
			mem[15] <=  32'b0_10000000_00000000000000000000000;  // 2;
			
			
			//	5.0: 	32'b01000000101000000000000000000000
			//	10.0: 	32'b01000001001000000000000000000000
			mem[16] <= 32'b01000100111110100000000000000000; //2000;
			mem[17] <= 32'b01000101000111000100000000000000; //2500;
			mem[18] <= 32'b01000101001110111000000000000000; //3000;
			mem[19] <= 32'b01000101010110101100000000000000; //3500;
			mem[20] <= 32'b01000101011110100000000000000000; //4000;
			mem[21] <= 32'b01000101100011001010000000000000; //4500;
			mem[22] <= 32'b01000101100111000100000000000000; //5000;
			mem[23] <= 32'b01000101101010111110000000000000; //5500;
			mem[24] <= 32'b01000101101110111000000000000000; //6000;
			mem[25] <= 32'b01000101110010110010000000000000; //6500;
			mem[26] <= 32'b01000101110110101100000000000000; //7000;
			mem[27] <= 32'b01000101111010100110000000000000; //7500;
			mem[28] <= 32'b01000101111110100000000000000000; //8000;
			mem[29] <= 32'b01000110000001001101000000000000; //8500;
			mem[30] <= 32'b01000110000011001010000000000000; //9000;
			mem[31] <= 32'b01000110000101000111000000000000; //9500;
			mem[32] <= 32'b01000110000111000100000000000000; //10000;
			mem[33] <= 32'b01000110001001000001000000000000; //10500;
			mem[34] <= 32'b01000110001010111110000000000000; //11000;
			mem[35] <= 32'b01000110001100111011000000000000; //11500;
			mem[36] <= 32'b01000110001110111000000000000000; //12000;
			mem[37] <= 32'b01000110010000110101000000000000; //12500;
			mem[38] <= 32'b01000110010010110010000000000000; //13000;
			mem[39] <= 32'b01000110010100101111000000000000; //13500;
			mem[40] <= 32'b01000110010110101100000000000000; //14000;
			mem[41] <= 32'b01000110011000101001000000000000; //14500;
			mem[42] <= 32'b01000110011010100110000000000000; //15000;
			mem[43] <= 32'b01000110011100100011000000000000; //15500;
			mem[44] <= 32'b01000110011110100000000000000000; //16000;
			mem[45] <= 32'b01000110100000001110100000000000; //16500;
			mem[46] <= 32'b01000110100001001101000000000000; //17000;
			mem[47] <= 32'b01000110100010001011100000000000; //17500;
			
			mem[64]  <=  32'b0_10000000_00000000000000000000000;  //2.0;
			mem[66]  <=  32'b0_10000001_00000000000000000000000;  //4.0;
			mem[68]  <=  32'b0_10000001_10000000000000000000000;  //6.0;
			mem[70]  <=  32'b0_10000010_00000000000000000000000;  //8.0;
			mem[72]  <=  32'b0_10000010_01000000000000000000000;  //10.0;
			mem[74]  <=  32'b0_10000010_10000000000000000000000;  //12.0;
			mem[76]  <=  32'b0_10000010_11000000000000000000000;  //14.0;
			mem[78]  <=  32'b0_10000011_00000000000000000000000;  //16.0;
			mem[80]  <=  32'b0_10000011_00100000000000000000000;  //18.0;
			mem[82]  <=  32'b0_10000011_01000000000000000000000;  //20.0;
			mem[84]  <=  32'b0_10000011_01100000000000000000000;  //22.0;
			mem[86]  <=  32'b0_10000011_10000000000000000000000;  //24.0;
			mem[88]  <=  32'b0_10000011_10100000000000000000000;  //26.0;
			mem[90]  <=  32'b0_10000011_11000000000000000000000;  //28.0;
			mem[92]  <=  32'b0_10000011_11100000000000000000000;  //30.0;
			mem[94]  <=  32'b0_10000100_00000000000000000000000;  //32.0;
			mem[96]  <=  32'b0_10000100_00010000000000000000000;  //34.0;
			mem[98]  <=  32'b0_10000100_00100000000000000000000;  //36.0;
			mem[100] <=  32'b0_10000100_00110000000000000000000;  //38.0;
			mem[102] <=  32'b0_10000100_01000000000000000000000;  //40.0;
			mem[104] <=  32'b0_10000100_01010000000000000000000;  //42.0;
			mem[106] <=  32'b0_10000100_01100000000000000000000;  //44.0;
			mem[108] <=  32'b0_10000100_01110000000000000000000;  //46.0;
			mem[110] <=  32'b0_10000100_10000000000000000000000;  //48.0;
			mem[112] <=  32'b0_10000100_10010000000000000000000;  //50.0;
			mem[114] <=  32'b0_10000100_10100000000000000000000;  //52.0;
			mem[116] <=  32'b0_10000100_10110000000000000000000;  //54.0;
			mem[118] <=  32'b0_10000100_11000000000000000000000;  //56.0;
			mem[120] <=  32'b0_10000100_11010000000000000000000;  //58.0;
			mem[122] <=  32'b0_10000100_11100000000000000000000;  //60.0;
			mem[124] <=  32'b0_10000100_11110000000000000000000;  //62.0;
			mem[126] <=  32'b0_10000101_00000000000000000000000;  //64.0;
    	end else if (w_en) begin
    		mem[addr_write] <= data;
    	end
    end
    
    // Bloque generate para asignar el espacio de rd_o a cada puerto
    // Parte baja al puerto 0
    // Parte alta al puerto 1
    generate
        genvar out;
        for (out = 0; out < MEM_READ_PORTS; out = out + 1) begin: mem_out_gen
            assign rd_o[out*WIDTH +: WIDTH] = mem[addr_read[out*DEPTH +: DEPTH]];
        end
    endgenerate
    
    
    // Bloque initial para asignar todos los contenidos de memoria a 0 nada más empezar
    initial begin
    	for(rst_mem = 0; rst_mem < 2**DEPTH; rst_mem = rst_mem + 1) begin
			mem[rst_mem] <= 0;
		end
    end
    
    // synthesis translate_on
  	
    reg [15:0] tics;
    always @(posedge clk) begin
    	if (rst) begin
    		tics <= 0;
    	end else begin
    		tics <= tics + 1;
    	end
    end
    
//    real float_aux = data;
    
    generate
        always @(posedge clk) begin
            if (w_en) begin
                $display ("Escritura memoria : posición %d : escrito = %.3f : ciclo %d", addr_write, data, tics);
            end
        end
    endgenerate
    // synthesis translate_on
    
endmodule
