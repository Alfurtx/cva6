// Original Author: Alfonso Amorós
// `include "vecunit/unit_dec_mem.sv"

module cvxif_unidad_vectorial_director
#(
) (
    input logic clk_i,
    input logic rst_i,
    input logic issue_valid
);

// Recibe una issue (comprobar issue_valid)
always_comb begin
end

endmodule
